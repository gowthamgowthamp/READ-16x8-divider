`include "Read_16x8.v"
`timescale 1ns/1ns
module Read_16x8_tb;
    reg [15:0]x;
    reg [7:0]y;
    reg bin;
    wire [7:0]q;
    wire [7:0]r;
    reg [7:0]app1;
    reg [7:0]app2;
    reg [7:0]app3;
    reg [7:0]app4;
    reg [7:0]app5;
    reg [7:0]app6;
    reg [7:0]app7;
    reg [7:0]app8;
    array error (.x(x), .y(y), .bin(bin), .q(q), .r(r), .app1(app1), .app2(app2), .app3(app3), .app4(app4), .app5(app5), .app6(app6), .app7(app7), .app8(app8));
    initial begin
        $dumpfile("Read_16x8_tb.vcd");
        $dumpvars(0, Read_16x8_tb);
        app1 = 255; app2 = 255; app3 = 255; app4 = 255; app5 = 255; app6 = 255; app7 = 255; app8 = 255; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 255; app3 = 255; app4 = 255; app5 = 255; app6 = 255; app7 = 254; app8 = 252; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 255; app3 = 255; app4 = 255; app5 = 255; app6 = 254; app7 = 252; app8 = 248; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 255; app3 = 255; app4 = 255; app5 = 254; app6 = 252; app7 = 248; app8 = 240; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 255; app3 = 255; app4 = 254; app5 = 252; app6 = 248; app7 = 240; app8 = 224; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 255; app3 = 254; app4 = 252; app5 = 248; app6 = 240; app7 = 224; app8 = 192; bin = 0;
                x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 255; app2 = 254; app3 = 252; app4 = 248; app5 = 240; app6 = 224; app7 = 192; app8 = 128; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
        app1 = 254; app2 = 252; app3 = 248; app4 = 240; app5 = 224; app6 = 192; app7 = 128; app8 = 0; bin = 0;
        x = 8; y = 4; #20;
        x = 7; y = 3; #20;
        x = 5; y = 5; #20;
        x = 16; y = 4; #20;
        x = 20; y = 5; #20;
        x = 15; y = 3; #20;
        x = 12; y = 5; #20;
        x = 40; y = 13; #20;
        x = 17; y = 5; #20;
        x = 199; y = 7; #20;
        x = 127; y = 5; #20;
    end
endmodule